* Rim et al. (2025) RLC Circuit - Step Response
* Tests transient response with step input at resonant frequency
*
* This validates the framework's ability to track envelope dynamics.

* ────────────────────────────────────────────────────────────
* PARAMETERS
* ────────────────────────────────────────────────────────────

.param Lval=100.04u
.param Cval=30.07n
.param Rs=3.0
.param Ro=2k
.param fres={1/(2*pi*sqrt(Lval*Cval))}

* ────────────────────────────────────────────────────────────
* CIRCUIT WITH STEP MODULATION
* ────────────────────────────────────────────────────────────

* Carrier source at resonant frequency
V1 N001 N002 SINE(0 1 {fres})

* Step modulation (0→1V at t=0.1ms)
Vmod N002 0 PULSE(0 1 0.1m 1n 1n 10m)

* Circuit
R1 N001 N003 {Rs}
L1 N003 N004 {Lval}
C1 N004 0 {Cval}
R2 N004 0 {Ro}

* ────────────────────────────────────────────────────────────
* SIMULATION
* ────────────────────────────────────────────────────────────

* Longer simulation to capture full transient
.tran 0 1m 0 1u

.save all

* Measure settling time
.meas TRAN Vfinal FIND V(N004) AT 1m
.meas TRAN Tsettle WHEN V(N004)=0.63*Vfinal RISE=1

.end
